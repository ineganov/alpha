`define HTRANS_IDLE    2'b00
`define HTRANS_NONSEQ  2'b10

`define HSIZE_1        3'b000
`define HSIZE_2        3'b001
`define HSIZE_4        3'b010
`define HSIZE_8        3'b011
